
interface intf(input logic clk,reset);
  
  //declaring the signals
  logic       valid;
  logic  a;
  logic  b;
  logic  c;
  logic  d;
  logic  out;
  logic  [1:0] sel;
  
endinterface